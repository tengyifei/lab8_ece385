module font_rom_32_bit ( input [10:0]	addr1,addr2,
						output [35:0]	data1, data2,
					 );

	parameter ADDR_WIDTH = 11;
   parameter DATA_WIDTH =  36;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
        
		  
36'b000000000000010010010000000000000000,
36'b000000000000000100100000000000000000,
36'b000000000000000101100000000000000000,
36'b000000000000101101101000000000000000,
36'b000000000000101100101000000000000000,
36'b000000000000101100101000000000000000,
36'b000000000000101100101000000000000000,
36'b000000000000010010010000000000000000,
36'b000000000000000010010000000000000000,
36'b000000000000000100100000000000000000,
36'b000000000000000100100000000000000000,
36'b000000000000000100100100000000000000
		  
		  
		  
		  
        };

	assign data1 = ROM[addr1];
	assign data2 = ROM[addr2];

endmodule  